
`include "defines.svh"
`include "des_if.svh"
`include "uvm_macros.svh"

package prj_pkg;
	import uvm_pkg::*;
	`include "uvm_sequence_item.svh"
	`include "uvm_monitor.svh"
	`include "uvm_scoreboard.svh"
	`include "uvm_driver.svh"
	`include "uvm_sequence.svh"
	`include "uvm_agent.svh"
	`include "uvm_env.svh"
	`include "uvm_test.svh"
endpackage
